../roms/characters.vh