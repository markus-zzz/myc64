../roms/basic.vh