../roms/kernal.vh